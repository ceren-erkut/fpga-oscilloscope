library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 
use IEEE.std_logic_unsigned.all; 
use ieee.numeric_std.ALL;

entity font_rom is Port (selectchar11: in integer; 
                         selectchar12: in integer; 
                         selectchar21: in integer; 
                         selectchar22: in integer; 
                         selectchar31: in integer; 
                         selectchar32: in integer; 
                         userlevel: in integer; 
                         mp1: in std_logic;mp2: in std_logic;
                         mp3: in std_logic;
                         display, Halfclock : in std_logic;
                         Rin, Bin, Gin : out std_logic_vector(3 downto 0);
                         pixel_X : in std_logic_vector(10 downto 0); 
                         pixel_Y : in std_logic_vector(9 downto 0); 
                         selectedY : in std_logic_vector(8 downto 0); 
                         selectedX: in std_logic_vector(9 downto 0));
end font_rom;
  
architecture Behavioral of font_rom is

type meas1 is array (0 to 32, 0 to 152) of std_logic; 
type meas2 is array (0 to 32, 0 to 152) of std_logic; 
type meas3 is array (0 to 32, 0 to 152) of std_logic; 
type char_rom2 is array (0 to 31, 0 to 15) of std_logic; 
type char_rom is array (0 to 15, 0 to 7) of std_logic;

constant vminString: meas3 := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0' ,'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1',' 1','1','0','0','1','1','0','0','1','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1 ','1','0','0 ','0','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0' ,'0','0','0','1',' 1','1','0','0','1','1','0','0','1','1','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','1','0','0','0 ','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','0','0','0','1','1',' 1','1','0','0','1','1','0','0','1','1','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1 ','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0',' 0','1','0',' 1','1','0','0','1','1','0','0','1','1','0','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','1 ','1','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','1','1','0',' 1','1','0','0','1','1','0','0','1','1','0','1','1','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','0 ','0','0','1 ','1','0','0','0','0','0','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','1','1','0','0','1','0','0','0','1','0','0','0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','0',' 1','1','0',' 1','1','0','0','1','1','0','0','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0', '1','1','1','0','0',' 1','1','0','0','1','1','0','0','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','0','0 ','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','1','1','1','1','1','1','1','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','1','0','0',' 1','1','0','0','1','1','0','0','1','1','0','0','0','1','1','1','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0 ','0','0','1 ','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','0','0' ,'0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1',' 0','0','0',' 1','1','0','0','1','1','0','0','1','1','0','0','0','1','1','1','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0 ','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','0','0','0','1','1','0','0','0','0','0','1','1','0' ,'0','0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1' ,'1','1','1', '0','0','1','1','1','1','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','0','0','0','1','1','0','0','0','0','1','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','1','1','0','0','1','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1' ,'0','0','0', '0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','1','1 ','0','0','0','0','1','1','0','0','1','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','0','1','1','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1' ,'0','0','0', '0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1' ,'0','0','0', '0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0', '0','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','1 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));                               
                    
constant vmaxString: meas2 :=(('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0' ,'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','1','1','1','0',' 0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1 ','1','0','0 ','0','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1', '1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1',' 1','1','0',' 0','0','0','1','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0 ','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','1','0','0','0','0' ,'0','1','1', '0','0','0','0','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','0','0','0','1','1','1','1','0',' 0','0','0','1','0','1','1','0','0','0','0','1','1','0','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1 ','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0' ,'0','1','0','0','0','0','0','0','1','0','1','1','0','0','0','1','1','0', '0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','0','0','0','1','0',' 1','1','0',' 0','0','1','1','0','1','1','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','1','1','0','0','0' ,'1','1','0', '0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','1','1','0',' 1','1','0',' 0','0','1','1','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','0 ','0','0','1 ','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','1',' 0','0','0','1','1','0', '0','1','1','1','1','0','0','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','0','1','1','0','1','1','0',' 0','1','1','0','0','0','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0 ','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0' , '0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','1','0','0',' 1','1','0',' 0','1','1','1','1','1','1','1','0','0','0','1','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','1','0','0','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','0','0' ,'1','1','0', '0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','1','1','0','0','1','1','1','0','0','1','1','0',' 0','1','0','0','0','0','0','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0 ','0','0','1 ','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1', '0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0',' 1','1','0',' 1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','0 ','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','0','0','0','1','1','0','0','0','0','0','1','1','0' ,'0','0','1', '1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' , '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1' ,'1','1','1', '0','0','1','1','1','1','0','0','1','1','0','0','0','0','0','0'),  
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','1','1','0','0','1','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0 ','0','0', '0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','1','1','0','0','1','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','0','1','1','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0',' 0','0','0','0','0','1','1','0','0', '0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0' ,'0','0','0','0','0','1','0','0','0', '0','1','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1' ,'1','0','0', '0','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));

constant vppString: meas1 := (('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','1','1','1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0', '1','1','0', '0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','1','1','0','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','1',' 1','1','1','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1 ','0','0','0 ','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','0','0','0','0','1','1', '1','1','1','0','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','1','1','0','0', '0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0',' 1','1','0',' 0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','0','0','0','1 ','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0','0','0' ,'1','1','0', '0','0','0','1','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','0','1','1','0','0','0','1','1','0','1','1', '0','0','0', '0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','1','1','0',' 0','0','0','0','0','0','1','0','1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','0 ','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','0','1','0','1','1','0','0','0','1','1','0','0', '0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','1','0','0','1','1','0','0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','1 ','1','0','0','0','0', '0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','1','1','0',' 1','1','0',' 0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1 ','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','0','1','0','0','0','0','0','1','1','0','1','1','0','0','0','1' ,'1','0','0', '0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','1','1','0','0','1','1','1','1','1','0','0','0','1','1','0','0','1','0','0','0','1','1','1','1','0','0','0','0', '0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0',' 1','1','1',' 1','1','0','0','0','1','0','0','0','1','1','0','0','1','1','1','1','0','0','0','0','0','0','0','0','1','1','0','0','1','0','0 ','0','1','1 ','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','0','0','0','1','1' ,'0','0','1','1','0','0', '1','1','1','1','0','0','1','1','1','1','1','0','0','0','0','0'),
('0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','1','1', '0','0','0', '0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0',' 0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','1','1','0','0 ','0','1','1 ','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0',' 0', '0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',' 0','0','1','1','1','1','1','1','1','0','0','1','1','0','1','1','1','0','0', '0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0',' 1','1','0',' 0','0','0','0','1','1','1','1','1','1','1','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','1','1','0','0','0','1','1 ','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','1','1','0','0','1' ,'1','0','0', '0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','1','1','0','0','1', '1','0','0', '0','0','0','0','0','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',' 0','0','0','0','1','0','0','0','0','0','1','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0','0','0 ','0','1','1 ','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0','0','1','0','0','0','0','0','1','1','0','0','1','1','0', '0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0'),
('0','0','1','1','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1','0','1','1' ,'0','0','0','1','1','0', '0','0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0',' 1','1','1',' 1','1','1','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0' ,'0','0','1','1','1','0','0','0','0','0','0 ','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','0' ,'0','1','1', '1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','1','1','1','1' ,'1','1','1', '0','0','1','1','1','1','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0 ','0','0','0','0','1','1','0','0', '0','1','1','0','0','1','0','0','0','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0' ,'0','0','0','0','0','1','1','0','0', '0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','0','1','1','0','0','1','0','0','0','1','1','0','0','0','0','0','1','0','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','0','1','1','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','0','0','0', '0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1 ','0','0','0','0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1' ,'1','0','0', '0','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','1','1','0','0', '0','1','0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','1','1 ','0','0','0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0','0','1','1','1','1','1','0','0','0','1' ,'1','0','0', '0','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1 ','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0' ,'0','0','0', '0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0', '0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0 ','0','0','0 ','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',' 0','0','0','0','0','0','0','0','0','0','0', '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));
  
constant number0 : char_rom2 :=( ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 3 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 3 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 4 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 4 
  ('1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0'), -- 5 
  ('1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0'), -- 5 
  ('1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0'), -- 6  
  ('1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0'), 
  ('1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','1','1','0','0','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'));

constant number1 : char_rom2 :=( ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 2 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 2 
  ('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'), -- 3 
  ('0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','0'), -- 3 
  ('0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0'), -- 4 
  ('0','0','1','1','1','1','1','1','1','1','0','0','0','0','0','0'), -- 4 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 5 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 5 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 6 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 6 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 7 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 7 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 8 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 8 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 9 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 9 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- a 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- a 
  ('0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0'), -- b 
  ('0','0','1','1','1','1','1','1','1','1','1','1','1','1','0','0'), -- b 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- d
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- e 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- d ****** 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- e 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')); -- f);

constant number2 : char_rom2 :=( ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 3 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 3 
  ('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0'), -- 4 
  ('0','0','0','0','0','0','0','0','0','0','1','1','1','1','0','0'), -- 4 
  ('0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0'), -- 5 
  ('0','0','0','0','0','0','0','0','1','1','1','1','0','0','0','0'), -- 5 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 6 
  ('0','0','0','0','0','0','1','1','1','1','0','0','0','0','0','0'), -- 6 
  ('0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0'), -- 7 
  ('0','0','0','0','1','1','1','1','0','0','0','0','0','0','0','0'), -- 7 
  ('0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'), -- 8 
  ('0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0'), -- 8 
  ('1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'), -- 9 
  ('1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0'), -- 9 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- a 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- a 
  ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'), -- b 
  ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0'), -- b 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- c 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')); -- f

constant number3 : char_rom2 :=( ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 0 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'), -- 1 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('0','0','1','1','1','1','1','1','1','1','1','1','0','0','0','0'), -- 2 
  ('1','1','1','1','0','0','0','0','0','0','1','1','1','1','0','0'), -- 3
  
  
  
  
  
  
  

